`timescale 1us/1ns

module MIPS_tb();

/////////////////////////////////////////////////////////
///////////////////// Parameters ////////////////////////
/////////////////////////////////////////////////////////
parameter CLK_PERIOD = 0.125 ;		//in us units


////////////////////////////////////////////////////////
/////////////////// DUT Signals //////////////////////// 
////////////////////////////////////////////////////////

reg					CLK_tb ;
reg					RST_tb ;
wire	[15:0] 		test_value_tb ;
////////////////////////////////////////////////////////
////////////////// initial block /////////////////////// 
////////////////////////////////////////////////////////
initial
 begin

  // Save Waveform
  $dumpfile("MIPS.vcd") ;       
  $dumpvars; 
  
  initialize();
  
  reset();
  


 #(100*CLK_PERIOD)
 $finish;
 end


////////////////////////////////////////////////////////
/////////////////////// TASKS //////////////////////////
////////////////////////////////////////////////////////
task initialize;
 begin
  CLK_tb = 1'b0;
 end
endtask 

task reset;
 begin
  RST_tb = 1'b1;
  #(CLK_PERIOD)
  RST_tb = 1'b0;
  #(CLK_PERIOD)
  RST_tb = 1'b1;
 end
endtask

////////////////////////////////////////////////////////
////////////////// Clock Generator  ////////////////////
////////////////////////////////////////////////////////
initial
 begin
	forever #(0.5*CLK_PERIOD)  CLK_tb = ~CLK_tb ;
 end
  
////////////////////////////////////////////////////////
/////////////////// DUT Instantation ///////////////////
////////////////////////////////////////////////////////
MIPS 	DUT(
.CLK(CLK_tb),
.RST(RST_tb),

.test_value(test_value_tb)
);



endmodule